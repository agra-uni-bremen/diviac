module divider_array_triangular_4_approx_div_49_57(n,d,q,r);
input [15:0]n;
input [7:0]d;
output [7:0]q,r;
 
wire [15:0]n1;
wire [7:0]d1;
wire [7:0]q1,r1;
wire [7:0]q,r;
wire [7:0]bout_local[0:7];
wire [7:0]r_local[0:7];
 
assign n1 = n;
assign d1 = d;
assign q = q1;
assign r = r1;
approx_div_49_57 sb0(n1[0],d1[0],1'b0,q1[0],r_local[0][0],bout_local[0][0]);
approx_div_49_57 sb1(n1[1],d1[0],1'b0,q1[1],r_local[1][0],bout_local[1][0]);
approx_div_49_57 sb2(n1[2],d1[0],1'b0,q1[2],r_local[2][0],bout_local[2][0]);
approx_div_49_57 sb3(n1[3],d1[0],1'b0,q1[3],r_local[3][0],bout_local[3][0]);
subtractor sb4(n1[4],d1[0],1'b0,q1[4],r_local[4][0],bout_local[4][0]);
subtractor sb5(n1[5],d1[0],1'b0,q1[5],r_local[5][0],bout_local[5][0]);
subtractor sb6(n1[6],d1[0],1'b0,q1[6],r_local[6][0],bout_local[6][0]);
subtractor sb7(n1[7],d1[0],1'b0,q1[7],r_local[7][0],bout_local[7][0]);
subtractor sb8(n1[8],d1[1],bout_local[7][0],q1[7],r_local[7][1],bout_local[7][1]);
subtractor sb9(n1[9],d1[2],bout_local[7][1],q1[7],r_local[7][2],bout_local[7][2]);
subtractor sb10(n1[10],d1[3],bout_local[7][2],q1[7],r_local[7][3],bout_local[7][3]);
subtractor sb11(n1[11],d1[4],bout_local[7][3],q1[7],r_local[7][4],bout_local[7][4]);
subtractor sb12(n1[12],d1[5],bout_local[7][4],q1[7],r_local[7][5],bout_local[7][5]);
subtractor sb13(n1[13],d1[6],bout_local[7][5],q1[7],r_local[7][6],bout_local[7][6]);
subtractor sb14(n1[14],d1[7],bout_local[7][6],q1[7],r_local[7][7],bout_local[7][7]);
approx_div_49_57 sb15(r_local[1][0],d1[1],bout_local[0][0],q1[0],r_local[0][1],bout_local[0][1]);
approx_div_49_57 sb16(r_local[1][1],d1[2],bout_local[0][1],q1[0],r_local[0][2],bout_local[0][2]);
approx_div_49_57 sb17(r_local[1][2],d1[3],bout_local[0][2],q1[0],r_local[0][3],bout_local[0][3]);
subtractor sb18(r_local[1][3],d1[4],bout_local[0][3],q1[0],r_local[0][4],bout_local[0][4]);
subtractor sb19(r_local[1][4],d1[5],bout_local[0][4],q1[0],r_local[0][5],bout_local[0][5]);
subtractor sb20(r_local[1][5],d1[6],bout_local[0][5],q1[0],r_local[0][6],bout_local[0][6]);
subtractor sb21(r_local[1][6],d1[7],bout_local[0][6],q1[0],r_local[0][7],bout_local[0][7]);
approx_div_49_57 sb22(r_local[2][0],d1[1],bout_local[1][0],q1[1],r_local[1][1],bout_local[1][1]);
approx_div_49_57 sb23(r_local[2][1],d1[2],bout_local[1][1],q1[1],r_local[1][2],bout_local[1][2]);
subtractor sb24(r_local[2][2],d1[3],bout_local[1][2],q1[1],r_local[1][3],bout_local[1][3]);
subtractor sb25(r_local[2][3],d1[4],bout_local[1][3],q1[1],r_local[1][4],bout_local[1][4]);
subtractor sb26(r_local[2][4],d1[5],bout_local[1][4],q1[1],r_local[1][5],bout_local[1][5]);
subtractor sb27(r_local[2][5],d1[6],bout_local[1][5],q1[1],r_local[1][6],bout_local[1][6]);
subtractor sb28(r_local[2][6],d1[7],bout_local[1][6],q1[1],r_local[1][7],bout_local[1][7]);
approx_div_49_57 sb29(r_local[3][0],d1[1],bout_local[2][0],q1[2],r_local[2][1],bout_local[2][1]);
subtractor sb30(r_local[3][1],d1[2],bout_local[2][1],q1[2],r_local[2][2],bout_local[2][2]);
subtractor sb31(r_local[3][2],d1[3],bout_local[2][2],q1[2],r_local[2][3],bout_local[2][3]);
subtractor sb32(r_local[3][3],d1[4],bout_local[2][3],q1[2],r_local[2][4],bout_local[2][4]);
subtractor sb33(r_local[3][4],d1[5],bout_local[2][4],q1[2],r_local[2][5],bout_local[2][5]);
subtractor sb34(r_local[3][5],d1[6],bout_local[2][5],q1[2],r_local[2][6],bout_local[2][6]);
subtractor sb35(r_local[3][6],d1[7],bout_local[2][6],q1[2],r_local[2][7],bout_local[2][7]);
subtractor sb36(r_local[4][0],d1[1],bout_local[3][0],q1[3],r_local[3][1],bout_local[3][1]);
subtractor sb37(r_local[4][1],d1[2],bout_local[3][1],q1[3],r_local[3][2],bout_local[3][2]);
subtractor sb38(r_local[4][2],d1[3],bout_local[3][2],q1[3],r_local[3][3],bout_local[3][3]);
subtractor sb39(r_local[4][3],d1[4],bout_local[3][3],q1[3],r_local[3][4],bout_local[3][4]);
subtractor sb40(r_local[4][4],d1[5],bout_local[3][4],q1[3],r_local[3][5],bout_local[3][5]);
subtractor sb41(r_local[4][5],d1[6],bout_local[3][5],q1[3],r_local[3][6],bout_local[3][6]);
subtractor sb42(r_local[4][6],d1[7],bout_local[3][6],q1[3],r_local[3][7],bout_local[3][7]);
subtractor sb43(r_local[5][0],d1[1],bout_local[4][0],q1[4],r_local[4][1],bout_local[4][1]);
subtractor sb44(r_local[5][1],d1[2],bout_local[4][1],q1[4],r_local[4][2],bout_local[4][2]);
subtractor sb45(r_local[5][2],d1[3],bout_local[4][2],q1[4],r_local[4][3],bout_local[4][3]);
subtractor sb46(r_local[5][3],d1[4],bout_local[4][3],q1[4],r_local[4][4],bout_local[4][4]);
subtractor sb47(r_local[5][4],d1[5],bout_local[4][4],q1[4],r_local[4][5],bout_local[4][5]);
subtractor sb48(r_local[5][5],d1[6],bout_local[4][5],q1[4],r_local[4][6],bout_local[4][6]);
subtractor sb49(r_local[5][6],d1[7],bout_local[4][6],q1[4],r_local[4][7],bout_local[4][7]);
subtractor sb50(r_local[6][0],d1[1],bout_local[5][0],q1[5],r_local[5][1],bout_local[5][1]);
subtractor sb51(r_local[6][1],d1[2],bout_local[5][1],q1[5],r_local[5][2],bout_local[5][2]);
subtractor sb52(r_local[6][2],d1[3],bout_local[5][2],q1[5],r_local[5][3],bout_local[5][3]);
subtractor sb53(r_local[6][3],d1[4],bout_local[5][3],q1[5],r_local[5][4],bout_local[5][4]);
subtractor sb54(r_local[6][4],d1[5],bout_local[5][4],q1[5],r_local[5][5],bout_local[5][5]);
subtractor sb55(r_local[6][5],d1[6],bout_local[5][5],q1[5],r_local[5][6],bout_local[5][6]);
subtractor sb56(r_local[6][6],d1[7],bout_local[5][6],q1[5],r_local[5][7],bout_local[5][7]);
subtractor sb57(r_local[7][0],d1[1],bout_local[6][0],q1[6],r_local[6][1],bout_local[6][1]);
subtractor sb58(r_local[7][1],d1[2],bout_local[6][1],q1[6],r_local[6][2],bout_local[6][2]);
subtractor sb59(r_local[7][2],d1[3],bout_local[6][2],q1[6],r_local[6][3],bout_local[6][3]);
subtractor sb60(r_local[7][3],d1[4],bout_local[6][3],q1[6],r_local[6][4],bout_local[6][4]);
subtractor sb61(r_local[7][4],d1[5],bout_local[6][4],q1[6],r_local[6][5],bout_local[6][5]);
subtractor sb62(r_local[7][5],d1[6],bout_local[6][5],q1[6],r_local[6][6],bout_local[6][6]);
subtractor sb63(r_local[7][6],d1[7],bout_local[6][6],q1[6],r_local[6][7],bout_local[6][7]);
assign q1[0] = (r_local[1][7])|(~bout_local[0][7]); 
assign q1[1] = (r_local[2][7])|(~bout_local[1][7]); 
assign q1[2] = (r_local[3][7])|(~bout_local[2][7]); 
assign q1[3] = (r_local[4][7])|(~bout_local[3][7]); 
assign q1[4] = (r_local[5][7])|(~bout_local[4][7]); 
assign q1[5] = (r_local[6][7])|(~bout_local[5][7]); 
assign q1[6] = (r_local[7][7])|(~bout_local[6][7]); 
assign q1[7] = (n1[15])|(~bout_local[7][7]); 
assign r1[0] = r_local[0][0]; 
assign r1[1] = r_local[0][1]; 
assign r1[2] = r_local[0][2]; 
assign r1[3] = r_local[0][3]; 
assign r1[4] = r_local[0][4]; 
assign r1[5] = r_local[0][5]; 
assign r1[6] = r_local[0][6]; 
assign r1[7] = r_local[0][7]; 
endmodule 
module subtractor(x_exact,y_exact,bin_exact,qs_exact,r_sub_exact,bout_exact); 
 
input x_exact,y_exact,bin_exact,qs_exact; 
output r_sub_exact,bout_exact; 
wire diff_exact; 
assign diff_exact = x_exact^y_exact^bin_exact; 
assign bout_exact = (~x_exact & y_exact)|((~(x_exact^y_exact)) & bin_exact); 
assign r_sub_exact = qs_exact?diff_exact:x_exact; 
endmodule
module approx_div_49_57(x, y, bin, qs, r_sub, bout);
input x, y, bin, qs;
output r_sub, bout;
wire diff; 
assign bout = 0 | (~x & y & ~bin) | (~x & y & bin) | (x & y & bin) ;
assign diff = 0 | (~x & y & ~bin) | (~x & y & bin) | (x & ~y & ~bin) | (x & y & bin) ;
assign r_sub = qs?diff:x ;
endmodule
